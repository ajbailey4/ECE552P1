module cpu(clk, rst_n, hlt, pc);
	
	input clk, rst_n;
	output hlt;
	output [15:0] pc;
	
	
endmodule